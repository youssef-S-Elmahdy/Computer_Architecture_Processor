
module Memory (input clk, input MemRead, input MemWrite, input [2:0] funct3, input [7:0] addr, input [31:0] data_in, output reg [31:0] data_out);
       
    reg [7:0] mem [0:255]; 
    always @ (posedge clk) begin
        if(MemWrite) begin
            case(funct3)
                3'b000: mem[addr] <= data_in[7:0]; // SB
                3'b001: begin // SH
                    mem[addr] <= data_in[7:0];
                    mem[addr+1] <= data_in[15:8];
                end
                3'b010: begin // SW
                    mem[addr] <= data_in[7:0];
                    mem[addr+1] <= data_in[15:8];
                    mem[addr+2] <= data_in[23:16];
                    mem[addr+3] <= data_in[31:24];
                end
                default: begin 
                    mem[addr] <= data_in[7:0];
                    mem[addr+1] <= data_in[15:8];
                    mem[addr+2] <= data_in[23:16];
                    mem[addr+3] <= data_in[31:24];
                end
            endcase 
        end
        else
            mem[addr] <= mem[addr];
    end 
    
    always @ (*) begin
        if(MemRead) begin
            case(funct3)
                3'b000: data_out = {{24{mem[addr][7]}}, mem[addr]}; // LB
                3'b001: data_out = {{16{mem[addr+1][7]}}, mem[addr+1], mem[addr]}; // LH
                3'b010: data_out = {mem[addr+3], mem[addr+2], mem[addr+1], mem[addr]}; // LW
                3'b100: data_out = {24'b0, mem[addr]}; // LBU
                3'b101: data_out = {16'b0, mem[addr+1], mem[addr]}; // LHU
                default: data_out = {mem[addr+3], mem[addr+2], mem[addr+1], mem[addr]}; // LW
            endcase 
        end
        else
            data_out = 32'b0;
    end 
    initial begin
//    test case 1
//        {mem[3], mem[2], mem[1], mem[0]} = 32'b11111111101100000000000010010011; //addi x1, x0, -5 
//        {mem[7], mem[6], mem[5], mem[4]} = 32'b00000000001100001010000100010011; //slti x2, x1, 3
//        {mem[11], mem[10], mem[9], mem[8]} = 32'b00000000001100001011000110010011; //sltiu x3, x1, 3
//        {mem[15], mem[14], mem[13], mem[12]} = 32'b00000001010000011100001000010011; //xori x4, x3, 20
//        {mem[19], mem[18], mem[17], mem[16]} = 32'b00000101010100100110001010010011; //ori x5, x4, 85
//        {mem[23], mem[22], mem[21], mem[20]} = 32'b11111110011100001111001100010011; //andi x6, x1, -25
//        {mem[27], mem[26], mem[25], mem[24]} = 32'b00000000010000010001001110010011; //slli x7, x2, 4
//        {mem[31], mem[30], mem[29], mem[28]} = 32'b00000000001000100101010000010011; //srli x8, x4, 2
//        {mem[35], mem[34], mem[33], mem[32]} = 32'b01000000001000110101010010010011; //srai x9, x6, 2

//test case 2
//{mem[3], mem[2], mem[1], mem[0]} = 32'b00000000000100000000001010010011; //addi x5, x0, 1 # x = 1
//{mem[7], mem[6], mem[5], mem[4]} = 32'b00000000000000000000001100010011; //addi x6, x0, 0 # i = 0
//{mem[11], mem[10], mem[9], mem[8]} = 32'b00000000011000000000001110010011; //addi x7, x0, 6 # y = 6
//{mem[15], mem[14], mem[13], mem[12]} = 32'b00000000011100101000101001100011; //beq x5, x7, endStore # i == y?

//{mem[19], mem[18], mem[17], mem[16]} = 32'b00000000010100110010000000100011; //sw x5, 0(x6)
//{mem[23], mem[22], mem[21], mem[20]} = 32'b00000000010000110000001100010011; //addi x6, x6, 4
//{mem[27], mem[26], mem[25], mem[24]} = 32'b00000000000100101000001010010011; //addi x5, x5, 1
//{mem[31], mem[30], mem[29], mem[28]} = 32'b11111110000000000000100011100011; //beq x0, x0, store # loop back

//{mem[35], mem[34], mem[33], mem[32]} = 32'b00000000000000000000001010010011; //addi x5, x0, 0 # i = 0
//{mem[39], mem[38], mem[37], mem[36]} = 32'b00000000000000000000001100010011; //addi x6, x0, 0 # *i

//{mem[43], mem[42], mem[41], mem[40]} = 32'b00000001000000000000001110010011; //addi x7, x0, 16 # *(4-i)
//{mem[47], mem[46], mem[45], mem[44]} = 32'b00000000001100000000111000010011; //addi x8, x0, 3 # x = 3
//{mem[51], mem[50], mem[49], mem[48]} = 32'b00000011110000101000001001100011; //beq x5, x8, endSwap # i == x?
//{mem[55], mem[54], mem[53], mem[52]} = 32'b00000000000000110010111010000011; //lw x9, 0(x6) # temp1 = mem[i]
//{mem[59], mem[58], mem[57], mem[56]} = 32'b00000000000000111010111100000011; //lw x10, 0(x7) # temp2 = mem[4-i]
//{mem[63], mem[62], mem[61], mem[60]} = 32'b00000001110100111010000000100011; //sw x9, 0(x7) # mem[4-i] = temp1
//{mem[67], mem[66], mem[65], mem[64]} = 32'b00000001111000110010000000100011; //sw x10, 0(x6) # mem[i] = temp2

//{mem[71], mem[70], mem[69], mem[68]} = 32'b00000000000100101000001010010011; //addi x5, x5, 1 # i++
//{mem[75], mem[74], mem[73], mem[72]} = 32'b00000000010000110000001100010011; //addi x6, x6, 4 # *(i+1)
//{mem[79], mem[78], mem[77], mem[76]} = 32'b11111111110000111000001110010011; //addi x7, x7, -4 # *(4-i-1)
//{mem[83], mem[82], mem[81], mem[80]} = 32'b11111110000000000000000011100011; //beq x0, x0, swap # loop back

//Test case 3
//    {mem[3], mem[2], mem[1], mem[0]} = 32'b00000000000000000100000010000011; // lbu x1, 0(x0) #x1 = 24
//    {mem[7], mem[6], mem[5], mem[4]} = 32'b00000000010000000001000100000011; // lh x2, 4(x0) #x2 = 2
//    {mem[11], mem[10], mem[9], mem[8]} = 32'b00000000100000000000000110000011; // lb x3, 8(x0) #x3 = -126
//    {mem[15], mem[14], mem[13], mem[12]} = 32'b00000000110000000101001000000011; // lhu x4, 12(x0) #x4 = 3
//    {mem[19], mem[18], mem[17], mem[16]} =32'b00000000001000001001001010110011; // sll x5, x1, x2 #x5 = 96
//    {mem[23], mem[22], mem[21], mem[20]} = 32'b00000000000100011010001100110011; // slt x6, x3, x1 #x6 = 1
//    {mem[27], mem[26], mem[25], mem[24]} = 32'b00000000000100011011001110110011; // sltu x7, x3, x1 #x7 = 0
//    {mem[31], mem[30], mem[29], mem[28]} = 32'b00000000010100110100010000110011; // xor x8, x6, x5 #x8 = 97
//    {mem[35], mem[34], mem[33], mem[32]} = 32'b00000000001000011101010010110011; // srl x9, x3, x2 #x9 = 1073741792 
//    {mem[39], mem[38], mem[37], mem[36]} = 32'b01000000001000011101010100110011; // sra x10,x3, x2 #x10 = -32 
    
    
//    {mem[43], mem[42], mem[41], mem [40]} = 32'b00000000000000000000000000011000; // 24
//    {mem[47], mem[46], mem[45], mem[44]} = 32'b00000000000000000000000000000010; // 2
//    {mem[51], mem[50], mem[49], mem[48]} = 32'b00000000000000000000000010000010; // 66
//    {mem[55], mem[54], mem[53], mem[52]} = 32'b00000000000000000000000000000011; // 3

//Test case 4
//    {mem[3], mem[2], mem[1], mem[0]} = 32'b000000000000_00000_010_00001_0000011; // lw x1, 0(x0) 
//    {mem[7], mem[6], mem[5], mem[4]} = 32'b0000000_00000_00001_110_00100_0110011; // or x4, x1, x0 
//    {mem[11], mem[10], mem[9], mem[8]} = 32'b0000000_00100_00000_010_01100_0100011; // sw x4, 12(x0)
    
    
//    {mem[15], mem[14], mem[13], mem[12]} = 32'd15;


//Test case 5
//    {mem[3], mem[2], mem[1], mem[0]} = 32'b00000000000000000010000010110111; // lui x1, 2
//    {mem[7], mem[6], mem[5], mem[4]} = 32'b00000000000000000101000100010111; // auipc x2, 5    
//    {mem[11], mem[10], mem[9], mem[8]} = 32'b00000000100000000000000111101111; // jal x3, 8
     
//    {mem[15], mem[14], mem[13], mem[12]} = 32'b00000000000100000000000001110011; // ebreak 
//    {mem[19], mem[18], mem[17], mem[16]} = 32'b00000000001000001001010001100011; // bne x1, x2, 8
    
//    {mem[23], mem[22], mem[21], mem[20]} = 32'b00000000000000000000000001110011; // ecall 
//    {mem[27], mem[26], mem[25], mem[24]} = 32'b11111100100000000000001000010011; // addi x4, x0, -56
//    {mem[31], mem[30], mem[29], mem[28]} = 32'b00000000001000001100010001100011; // blt x1, x2, 8 
    
//    {mem[35], mem[34], mem[33], mem[32]} = 32'b00000000000000000000000001110011; // ecall 
//    {mem[39], mem[38], mem[37], mem[36]} = 32'b00000000001000000000000000100011; // sb x2, 0(x0) 
//    {mem[43], mem[42], mem[41], mem[40]} = 32'b00000000000100010101010001100011; // bge x2, x1, 8 
    
//    {mem[47], mem[46], mem[45], mem[44]} = 32'b00000000000000000000000001110011; // ecall
//    {mem[51], mem[50], mem[49], mem[48]} = 32'b00000000010000001110010001100011; // bltu x1, x4, 8 
    
//    {mem[55], mem[54], mem[53], mem[52]} = 32'b00000000000000000000000001110011; // ecall 
//    {mem[59], mem[58], mem[57], mem[56]} = 32'b00000000001000100111010001100011; // bgeu x4, x2, 8
      
//    {mem[63], mem[62], mem[61], mem[60]} = 32'b00000000000000000000000001110011; // ecall  
//    {mem[67], mem[66], mem[65], mem[64]} = 32'b00000000010000000001000010100011; // sh x4, 1(x0) 
//    {mem[71], mem[70], mem[69], mem[68]} = 32'b00000000000000000000000001110011; // ecall 
//    {mem[75], mem[74], mem[73], mem[72]} = 32'b00001111111100000000000000001111; // fence
//    {mem[79], mem[78], mem[77], mem[76]} = 32'b00000000000000011000000001100111; //  jalr x0, x3, 0

//Test case 6
//    {mem[3], mem[2], mem[1], mem[0]} = 32'b00000000000000000010000100000011; // lw x2, 0(x0)
//    {mem[7], mem[6], mem[5], mem[4]} = 32'b00000000010000000010000110000011; // lw x3, 4(x0)   
//    {mem[11], mem[10], mem[9], mem[8]} = 32'b00000000001100010000001000110011; // add x4, x2, x3
//    {mem[15], mem[14], mem[13], mem[12]} = 32'b01000000001100100000001010110011; // sub x5, x4, x3
//    {mem[19], mem[18], mem[17], mem[16]} = 32'b00000000001100010111001100110011; // and x6, x2, x3
    
//    {mem[23], mem[22], mem[21], mem[20]} = 32'b00000000000000000000000000000011; // 3 
//    {mem[27], mem[26], mem[25], mem[24]} = 32'b00000000000000000000000000000111; // 7
    end

endmodule 