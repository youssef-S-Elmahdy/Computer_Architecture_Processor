

module InstMem (input [5:0] addr, output [31:0] data_out); 
    reg [31:0] mem [0:63]; 
     
    initial begin 
        mem[0] = 32'b00000000100000001000000100010011; //addi x2,x1,8
        mem[1] = 32'b00000000000000010000000110110011; //add x3, x2, x0
        mem[2] = 32'b00000000000000001010001000000011; //lw x4,0(x1)
        mem[3] = 32'b00000000010000000010011000100011; //sw x4, 12(x0)
        mem[4] = 32'b00000000000000010000011001100011; //beq x2, x0, 12 "False"
        mem[5] = 32'b00000000001000011111001010110011; //and x5, x3, x2
        mem[6] = 32'b00000000000000101110010010110011; //or x9, x5, x0
        mem[7] = 32'b00000000000000001000010001100011; //beq x1,x0,8
        mem[8] = 32'b01000000000100010000000000110011; //sub x0, x2, x1
        mem[9] = 32'b00000000001000010001010000010011; //slli x8, x2, 2
        mem[10] = 32'b00000001100000000000000011101111; //jal x1, 24
        mem[16] = 32'b00000000001111101000011110110111; //lui x15, 1000
        mem[17] = 32'b00000000000001100100101000010111; //auipc x20, 100
        mem[18] = 32'b01000000111110100000101010110011; //sub x21, x20, x15
        mem[19] = 32'b00000000111100000110010001100011; //bltu x0, x15, 8
        mem[20] = 32'b00000000000000000000000010110011; //add x1, x0, x0
        mem[21] = 32'b00000000111110100010101100110011; //slt x22, x20, x15
        mem[22] = 32'b00000000010000000001010001100011; //bne x0, x4, 8
        mem[24] = 32'b00000000000000000001011001100011; //bne x0,x0,12 "False"
        mem[25] = 32'b11111111111111111111010100110111; //lui x10,1048575
        mem[26] = 32'b00000000010001010101010110010011; //srli x11, x10, 4
        mem[27] = 32'b01000000010001010101011000010011; //srai x12, x10, 4
        mem[28] = 32'b00000000000000011100001110010011; //xori x7, x3, 0
        mem[29] = 32'b00000000101000011011010000010011; //sltiu x8, x3, 10
        mem[30] = 32'b00000000000001111000000001100111; //jalr x0, 0(x15)
    end 
     
    assign data_out = mem[addr];
endmodule


